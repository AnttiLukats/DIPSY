library work;


package config is

	constant CFG_VENDOR : string := "sbt";
	constant CFG_BOARD : string := "st32ice";

	constant CFG_FIRST_IO : integer := 0;
	constant CFG_LAST_IO : integer := 4;


end;